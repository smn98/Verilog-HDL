`timescale 1ns / 1ps

module bin2ex3(
    input [2:0] b,
    output [3:0] e
    );

assign e = b + 3;

endmodule
